
module clock_gater(
    //--------------------------------------------------------------------------
    // Global signals
    //--------------------------------------------------------------------------
    clk,
    reset,

    //--------------------------------------------------------------------------
    // Input interface
    //--------------------------------------------------------------------------
    i__enable,

    //--------------------------------------------------------------------------
    // Output interface
    //--------------------------------------------------------------------------
    o__gated_clk
);

//------------------------------------------------------------------------------
// Global signals
//------------------------------------------------------------------------------
input  logic                            clk;
input  logic                            reset;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Iuput interface
//------------------------------------------------------------------------------
input  logic                            i__enable;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Output interface
//------------------------------------------------------------------------------
output logic                            o__gated_clk;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Signals
//------------------------------------------------------------------------------
logic                                   w__enable_latched;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Generate gated clock
//------------------------------------------------------------------------------
`ifndef USE_STDCELL_LATCH
always_latch
begin
    if(clk == 1'b0)
    begin
        w__enable_latched <= i__enable;
    end
end

always_comb
begin
    o__gated_clk = clk & w__enable_latched;
end
`else
//PREICG_X1B_A12TH
//    latch (
//        .CK                             (clk),
//        .SE                             (reset),
//        .E                              (i__enable),
//        .ECK                            (o__gated_clk)
//    );
`endif
//------------------------------------------------------------------------------

endmodule

