// `ifndef _pifo_incl_vh_ 
// `define _pifo_incl_vh_

import PifoPkg::*;

// `endif
