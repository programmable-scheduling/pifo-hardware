// `ifndef _pifo_tb_incl_vh_ 
// `define _pifo_tb_incl_vh_
import PifoTbPkg::*;

// `endif
