
module counter(
    //--------------------------------------------------------------------------
    // Global signals
    //--------------------------------------------------------------------------
    clk,
    reset,

    //--------------------------------------------------------------------------
    // Input interface
    //--------------------------------------------------------------------------
    i__inc,

    //--------------------------------------------------------------------------
    // Output interface
    //--------------------------------------------------------------------------
    o__count,
    o__count__next
);

//------------------------------------------------------------------------------
// Parameters
//------------------------------------------------------------------------------
parameter NUM_COUNT                     = 8;
parameter COUNT_WIDTH                   = $clog2(NUM_COUNT);
parameter INIT_VALUE                    = 1'b0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Global signals
//------------------------------------------------------------------------------
input  logic                            clk;
input  logic                            reset;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Input interface
//------------------------------------------------------------------------------
input  logic                            i__inc;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Output interface
//------------------------------------------------------------------------------
output logic [COUNT_WIDTH-1:0]          o__count;
output logic [COUNT_WIDTH-1:0]          o__count__next;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Internal signals
//------------------------------------------------------------------------------
logic [COUNT_WIDTH-1:0]                 w__max_count;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Submodules
//------------------------------------------------------------------------------
counter_base
    #(
        .COUNT_WIDTH                    (COUNT_WIDTH),
        .INIT_VALUE                     (INIT_VALUE)
    )
    base(
        .clk                            (clk),
        .reset                          (reset),
        .i__max_count                   (w__max_count),
        .i__inc                         (i__inc),
        .o__count                       (o__count),
        .o__count__next                 (o__count__next)
    );
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Max count logic
//------------------------------------------------------------------------------
always_comb
begin
    // To eliminate the 32-bit to ?-bit conversion warnings
    w__max_count = NUM_COUNT - 1'b1;
end
//------------------------------------------------------------------------------

endmodule

