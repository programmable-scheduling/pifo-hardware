// `ifndef _flow_pifo_tb_incl_vh_ 
// `define _flow_pifo_tb_incl_vh_
import FlowPifoTbPkg::*;
import InterfacePkg::*;
import CommonTbPkg::*;
import FlowPifoPkg::*;

// `endif
