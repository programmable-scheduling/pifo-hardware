// `ifndef _common_tb_incl_vh_ 
// `define _common_tb_incl_vh_
import CommonTbPkg::*;

// `endif
