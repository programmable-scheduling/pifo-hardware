module counter(
    //--------------------------------------------------------------------------
    // Global signals
    //--------------------------------------------------------------------------
    clk,
    reset,

    //--------------------------------------------------------------------------
    // Input interface
    //--------------------------------------------------------------------------
    i__inc,

    //--------------------------------------------------------------------------
    // Output interface
    //--------------------------------------------------------------------------
    o__count,
    o__count__next
);

//------------------------------------------------------------------------------
// Parameters
//------------------------------------------------------------------------------
parameter NUM_COUNT                     = 8;
parameter COUNT_WIDTH                   = $clog2(NUM_COUNT);
parameter INIT_VALUE                    = 1'b0;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Global signals
//------------------------------------------------------------------------------
input  logic                            clk;
input  logic                            reset;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Input interface
//------------------------------------------------------------------------------
input  logic                            i__inc;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Output interface
//------------------------------------------------------------------------------
output logic [COUNT_WIDTH-1:0]          o__count;
output logic [COUNT_WIDTH-1:0]          o__count__next;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Internal signals
//------------------------------------------------------------------------------
logic [COUNT_WIDTH-1:0]                 w__max_count;
logic [COUNT_WIDTH-1:0]                 r__count__pff;
logic [COUNT_WIDTH-1:0]                 w__count__next;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Output assignments
//------------------------------------------------------------------------------
assign o__count         = r__count__pff;
assign o__count__next   = w__count__next;
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Max count logic
//------------------------------------------------------------------------------
always_comb
begin
    // To eliminate the 32-bit to ?-bit conversion warnings
    w__max_count = NUM_COUNT - 1'b1;
end
//------------------------------------------------------------------------------

//------------------------------------------------------------------------------
// Count logic
//------------------------------------------------------------------------------
always_comb
begin
    w__count__next = r__count__pff;

    if(i__inc == 1'b1)
    begin
        if(r__count__pff == w__max_count)
        begin
            w__count__next = '0;
        end
        else
        begin
            w__count__next = r__count__pff + 1'b1;
        end
    end
end

always_ff @ (posedge clk)
begin
    if(reset == 1'b1)
    begin
        r__count__pff <= INIT_VALUE;
    end
    else
    begin
        r__count__pff <= w__count__next;
    end
end
//------------------------------------------------------------------------------

endmodule

